--------------------------------------------------------------------------------
-- nand_dumper_top.vhd
-- Top-level entity for the Arty Z7 NAND recovery design
--
-- This instantiates the AXI NAND controller and connects the NAND bus signals
-- to Pmod JA (data bus) and Pmod JB (control signals) through IOBUFs.
--
-- Pmod Pin Mapping:
--   JA[7:0]  -> NAND I/O[7:0]  (bidirectional data bus)
--   JB[0]    -> NAND CLE        (output)
--   JB[1]    -> NAND ALE        (output)
--   JB[2]    -> NAND CE#        (output, directly active low)
--   JB[3]    -> NAND WE#        (output, directly active low)
--   JB[4]    -> NAND RE#        (output, directly active low)
--   JB[5]    -> NAND WP#        (output, directly active low)
--   JB[6]    -> NAND R/B#       (input, directly active low)
--   JB[7]    -> spare / active-high LED for debug
--
-- Physical wiring: The desoldered NAND flash die must be connected to the
-- Pmod connectors via a breakout board or probe adapter. The NAND die pinout
-- must be identified first (typically from the die markings + ONFI datasheet).
--
-- Build flow: Use the Vivado Tcl script (tcl/create_project.tcl) to generate
-- the block design with the Zynq PS, then synthesize and implement.
--------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library unisim;
use unisim.vcomponents.all;

entity nand_dumper_top is
    port (
        -- Pmod JA: NAND data bus (directly to top-level bidirectional pads)
        JA : inout std_logic_vector(7 downto 0);

        -- Pmod JB: NAND control signals
        JB : inout std_logic_vector(7 downto 0);

        -- Fixed I/O for Zynq PS (directly to processing_system7 wrapper)
        DDR_addr          : inout std_logic_vector(14 downto 0);
        DDR_ba            : inout std_logic_vector(2 downto 0);
        DDR_cas_n         : inout std_logic;
        DDR_ck_n          : inout std_logic;
        DDR_ck_p          : inout std_logic;
        DDR_cke           : inout std_logic;
        DDR_cs_n          : inout std_logic;
        DDR_dm            : inout std_logic_vector(3 downto 0);
        DDR_dq            : inout std_logic_vector(31 downto 0);
        DDR_dqs_n         : inout std_logic_vector(3 downto 0);
        DDR_dqs_p         : inout std_logic_vector(3 downto 0);
        DDR_odt           : inout std_logic;
        DDR_ras_n         : inout std_logic;
        DDR_reset_n       : inout std_logic;
        DDR_we_n          : inout std_logic;
        FIXED_IO_ddr_vrn  : inout std_logic;
        FIXED_IO_ddr_vrp  : inout std_logic;
        FIXED_IO_mio      : inout std_logic_vector(53 downto 0);
        FIXED_IO_ps_clk   : inout std_logic;
        FIXED_IO_ps_porb  : inout std_logic;
        FIXED_IO_ps_srstb : inout std_logic
    );
end entity nand_dumper_top;

architecture structural of nand_dumper_top is

    ---------------------------------------------------------------------------
    -- Zynq PS wrapper component (generated by Vivado block design)
    -- The actual wrapper will be auto-generated. This declaration matches
    -- the standard Vivado PS7 wrapper with one M_AXI_GP0 port.
    ---------------------------------------------------------------------------
    component zynq_ps_wrapper is
        port (
            DDR_addr          : inout std_logic_vector(14 downto 0);
            DDR_ba            : inout std_logic_vector(2 downto 0);
            DDR_cas_n         : inout std_logic;
            DDR_ck_n          : inout std_logic;
            DDR_ck_p          : inout std_logic;
            DDR_cke           : inout std_logic;
            DDR_cs_n          : inout std_logic;
            DDR_dm            : inout std_logic_vector(3 downto 0);
            DDR_dq            : inout std_logic_vector(31 downto 0);
            DDR_dqs_n         : inout std_logic_vector(3 downto 0);
            DDR_dqs_p         : inout std_logic_vector(3 downto 0);
            DDR_odt           : inout std_logic;
            DDR_ras_n         : inout std_logic;
            DDR_reset_n       : inout std_logic;
            DDR_we_n          : inout std_logic;
            FIXED_IO_ddr_vrn  : inout std_logic;
            FIXED_IO_ddr_vrp  : inout std_logic;
            FIXED_IO_mio      : inout std_logic_vector(53 downto 0);
            FIXED_IO_ps_clk   : inout std_logic;
            FIXED_IO_ps_porb  : inout std_logic;
            FIXED_IO_ps_srstb : inout std_logic;
            -- FCLK
            FCLK_CLK0         : out std_logic;
            FCLK_RESET0_N     : out std_logic;
            -- M_AXI_GP0 (master from PS perspective, slave from PL perspective)
            M_AXI_GP0_ACLK    : in  std_logic;
            M_AXI_GP0_AWADDR  : out std_logic_vector(31 downto 0);
            M_AXI_GP0_AWVALID : out std_logic;
            M_AXI_GP0_AWREADY : in  std_logic;
            M_AXI_GP0_WDATA   : out std_logic_vector(31 downto 0);
            M_AXI_GP0_WSTRB   : out std_logic_vector(3 downto 0);
            M_AXI_GP0_WVALID  : out std_logic;
            M_AXI_GP0_WREADY  : in  std_logic;
            M_AXI_GP0_BRESP   : in  std_logic_vector(1 downto 0);
            M_AXI_GP0_BVALID  : in  std_logic;
            M_AXI_GP0_BREADY  : out std_logic;
            M_AXI_GP0_ARADDR  : out std_logic_vector(31 downto 0);
            M_AXI_GP0_ARVALID : out std_logic;
            M_AXI_GP0_ARREADY : in  std_logic;
            M_AXI_GP0_RDATA   : in  std_logic_vector(31 downto 0);
            M_AXI_GP0_RRESP   : in  std_logic_vector(1 downto 0);
            M_AXI_GP0_RVALID  : in  std_logic;
            M_AXI_GP0_RREADY  : out std_logic
        );
    end component;

    -- Clocks and resets from PS
    signal fclk_clk0    : std_logic;
    signal fclk_rstn    : std_logic;

    -- AXI GP0 signals
    signal gp0_awaddr   : std_logic_vector(31 downto 0);
    signal gp0_awvalid  : std_logic;
    signal gp0_awready  : std_logic;
    signal gp0_wdata    : std_logic_vector(31 downto 0);
    signal gp0_wstrb    : std_logic_vector(3 downto 0);
    signal gp0_wvalid   : std_logic;
    signal gp0_wready   : std_logic;
    signal gp0_bresp    : std_logic_vector(1 downto 0);
    signal gp0_bvalid   : std_logic;
    signal gp0_bready   : std_logic;
    signal gp0_araddr   : std_logic_vector(31 downto 0);
    signal gp0_arvalid  : std_logic;
    signal gp0_arready  : std_logic;
    signal gp0_rdata    : std_logic_vector(31 downto 0);
    signal gp0_rresp    : std_logic_vector(1 downto 0);
    signal gp0_rvalid   : std_logic;
    signal gp0_rready   : std_logic;

    -- NAND interface internal signals
    signal nand_io_i    : std_logic_vector(7 downto 0);
    signal nand_io_o    : std_logic_vector(7 downto 0);
    signal nand_io_t    : std_logic;
    signal nand_cle_i   : std_logic;
    signal nand_ale_i   : std_logic;
    signal nand_ce_n_i  : std_logic;
    signal nand_we_n_i  : std_logic;
    signal nand_re_n_i  : std_logic;
    signal nand_wp_n_i  : std_logic;
    signal nand_rb_n_i  : std_logic;

begin

    ---------------------------------------------------------------------------
    -- Zynq Processing System
    ---------------------------------------------------------------------------
    u_ps : zynq_ps_wrapper
        port map (
            DDR_addr          => DDR_addr,
            DDR_ba            => DDR_ba,
            DDR_cas_n         => DDR_cas_n,
            DDR_ck_n          => DDR_ck_n,
            DDR_ck_p          => DDR_ck_p,
            DDR_cke           => DDR_cke,
            DDR_cs_n          => DDR_cs_n,
            DDR_dm            => DDR_dm,
            DDR_dq            => DDR_dq,
            DDR_dqs_n         => DDR_dqs_n,
            DDR_dqs_p         => DDR_dqs_p,
            DDR_odt           => DDR_odt,
            DDR_ras_n         => DDR_ras_n,
            DDR_reset_n       => DDR_reset_n,
            DDR_we_n          => DDR_we_n,
            FIXED_IO_ddr_vrn  => FIXED_IO_ddr_vrn,
            FIXED_IO_ddr_vrp  => FIXED_IO_ddr_vrp,
            FIXED_IO_mio      => FIXED_IO_mio,
            FIXED_IO_ps_clk   => FIXED_IO_ps_clk,
            FIXED_IO_ps_porb  => FIXED_IO_ps_porb,
            FIXED_IO_ps_srstb => FIXED_IO_ps_srstb,
            FCLK_CLK0         => fclk_clk0,
            FCLK_RESET0_N     => fclk_rstn,
            M_AXI_GP0_ACLK    => fclk_clk0,
            M_AXI_GP0_AWADDR  => gp0_awaddr,
            M_AXI_GP0_AWVALID => gp0_awvalid,
            M_AXI_GP0_AWREADY => gp0_awready,
            M_AXI_GP0_WDATA   => gp0_wdata,
            M_AXI_GP0_WSTRB   => gp0_wstrb,
            M_AXI_GP0_WVALID  => gp0_wvalid,
            M_AXI_GP0_WREADY  => gp0_wready,
            M_AXI_GP0_BRESP   => gp0_bresp,
            M_AXI_GP0_BVALID  => gp0_bvalid,
            M_AXI_GP0_BREADY  => gp0_bready,
            M_AXI_GP0_ARADDR  => gp0_araddr,
            M_AXI_GP0_ARVALID => gp0_arvalid,
            M_AXI_GP0_ARREADY => gp0_arready,
            M_AXI_GP0_RDATA   => gp0_rdata,
            M_AXI_GP0_RRESP   => gp0_rresp,
            M_AXI_GP0_RVALID  => gp0_rvalid,
            M_AXI_GP0_RREADY  => gp0_rready
        );

    ---------------------------------------------------------------------------
    -- AXI NAND Controller
    -- PS GP0 AXI base address is typically 0x4000_0000.
    -- The lower 16 bits of the address are used for register/buffer access.
    ---------------------------------------------------------------------------
    u_axi_nand : entity work.axi_nand_ctrl
        generic map (
            C_S_AXI_DATA_WIDTH => 32,
            C_S_AXI_ADDR_WIDTH => 16,
            PAGE_BUF_DEPTH     => 18432
        )
        port map (
            s_axi_aclk    => fclk_clk0,
            s_axi_aresetn => fclk_rstn,
            s_axi_awaddr  => gp0_awaddr(15 downto 0),
            s_axi_awvalid => gp0_awvalid,
            s_axi_awready => gp0_awready,
            s_axi_wdata   => gp0_wdata,
            s_axi_wstrb   => gp0_wstrb,
            s_axi_wvalid  => gp0_wvalid,
            s_axi_wready  => gp0_wready,
            s_axi_bresp   => gp0_bresp,
            s_axi_bvalid  => gp0_bvalid,
            s_axi_bready  => gp0_bready,
            s_axi_araddr  => gp0_araddr(15 downto 0),
            s_axi_arvalid => gp0_arvalid,
            s_axi_arready => gp0_arready,
            s_axi_rdata   => gp0_rdata,
            s_axi_rresp   => gp0_rresp,
            s_axi_rvalid  => gp0_rvalid,
            s_axi_rready  => gp0_rready,
            nand_io_i     => nand_io_i,
            nand_io_o     => nand_io_o,
            nand_io_t     => nand_io_t,
            nand_cle      => nand_cle_i,
            nand_ale      => nand_ale_i,
            nand_ce_n     => nand_ce_n_i,
            nand_we_n     => nand_we_n_i,
            nand_re_n     => nand_re_n_i,
            nand_wp_n     => nand_wp_n_i,
            nand_rb_n     => nand_rb_n_i
        );

    ---------------------------------------------------------------------------
    -- Pmod JA: Bidirectional NAND data bus via IOBUFs
    ---------------------------------------------------------------------------
    gen_iobuf : for i in 0 to 7 generate
        u_iobuf : IOBUF
            generic map (
                DRIVE      => 12,
                IOSTANDARD => "DEFAULT",
                SLEW       => "SLOW"
            )
            port map (
                O  => nand_io_i(i),    -- FPGA input (from pad)
                IO => JA(i),           -- bidirectional pad
                I  => nand_io_o(i),    -- FPGA output (to pad)
                T  => nand_io_t        -- tristate: '1'=input, '0'=drive
            );
    end generate;

    ---------------------------------------------------------------------------
    -- Pmod JB: NAND control signals (directly driven outputs + R/B# input)
    ---------------------------------------------------------------------------
    JB(0) <= nand_cle_i;
    JB(1) <= nand_ale_i;
    JB(2) <= nand_ce_n_i;
    JB(3) <= nand_we_n_i;
    JB(4) <= nand_re_n_i;
    JB(5) <= nand_wp_n_i;

    -- R/B# is an input from the NAND (active low, open-drain)
    nand_rb_n_i <= JB(6);

    -- JB(7): debug output — directly mirror CE# for oscilloscope probing
    JB(7) <= nand_ce_n_i;

end architecture structural;
